`ifndef __TEST_WOR_V__
`define __TEST_WOR_V__

module test_wor(
	output wor y,
	input a, b, c, d, e, f, g, h, i
	);

	assign y = a;
	assign y = b;
	assign y = c;
	assign y = d;
	assign y = e;
	assign y = f;
	assign y = g;
	assign y = h;
	assign y = i;

endmodule

`endif /* __TEST_WOR_V__ */