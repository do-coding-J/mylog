.include lmv324.lib  ; LMV324 모델 라이브러리 파일 경로
* 모터 전류 회로

* 회로 정의
Vin in 0 DC 0V PULSE(0V 12V 0 1us 1us 1us 10ms)
R1 in 1 1k
XOPAMP 1 2 3 4 lmv324
R2 3 out 4.7k
C1 out 0 10n

* 시뮬레이션 설정
.tran 1us 10ms
.plot tran V(out)
.end
