* 네트리스트(회로) 정의
R1 1 0 1k       ; 1k 옴 저항
C1 1 2 10u      ; 10 마이크로 파라드 커패시터
V1 0 3 DC 5V    ; 5 볼트 DC 전원 공급

* 시뮬레이션 명령
.tran 1ms 10ms 0ms 1ms   ; 전이 응답 분석
.plot tran v(1) v(2)     ; 전압 v(1) 및 v(2) 그래프 플롯
.end