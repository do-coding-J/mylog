* LMV324 모델
* 모델 파라미터
.model LMV324 OPAMP (DC_GAIN=100K GBW=1M OFFSET=1mV CMRR=90dB)

* 회로 정의
Vin+ 1 0 DC 0V
Vin- 2 0 DC 0V
Vcc+ 7 0 DC 5V
Vcc- 8 0 DC -5V
Vout 6 0 DC 0V

* LMV324 Op-Amp 컴포넌트 정의
XOPAMP 1 2 6 LMV324

* 입력 신호 설정
V1 Vin+ 0 DC 1V
V2 Vin- 0 DC 0V

* 시뮬레이션 설정
.AC DEC 10 10Hz 100kHz
.TRAN 1ms 10ms

* 출력 플롯 설정
.plot AC Vdb(6)
.plot TRAN V(6)

* 시뮬레이션 실행
.AC Analysis
.TRAN Analysis
