VS N0 N1 DC 5V
R1 N1 N2 1K
C1 N2 0 1uF

.tran 1ms 10ms